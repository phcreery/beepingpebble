module fbg

import time
